* E:\Pr�ctica_3\Fuente_AC_RL_Vpulse.sch

* Schematics Version 9.1 - Web Update 1
* Thu May 18 09:56:19 2023



** Analysis setup **
.ac DEC 101 100 1000K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Fuente_AC_RL_Vpulse.net"
.INC "Fuente_AC_RL_Vpulse.als"


.probe


.END
