* E:\Pr�ctica_3\Fuente_AC_RC_Vpulse.sch

* Schematics Version 9.1 - Web Update 1
* Thu May 18 09:44:22 2023



** Analysis setup **
.tran 0.1ms 20ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Fuente_AC_RC_Vpulse.net"
.INC "Fuente_AC_RC_Vpulse.als"


.probe


.END
