* E:\Pr�ctica_3\Fuente_AC_RC.sch

* Schematics Version 9.1 - Web Update 1
* Thu May 18 10:03:41 2023



** Analysis setup **
.ac DEC 101 100 1000K
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Fuente_AC_RC.net"
.INC "Fuente_AC_RC.als"


.probe


.END
